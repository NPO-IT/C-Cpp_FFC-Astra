del_inst : del PORT MAP(
		clock	 => clock_sig,
		q	 => q_sig,
		cout	 => cout_sig
	);
