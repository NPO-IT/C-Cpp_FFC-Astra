count3_inst : count3 PORT MAP(
		clock	 => clock_sig,
		clk_en	 => clk_en_sig,
		q	 => q_sig,
		cout	 => cout_sig
	);
