compare_inst : compare PORT MAP(
		dataa	 => dataa_sig,
		AeB	 => AeB_sig
	);
