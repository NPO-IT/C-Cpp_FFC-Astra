compare4_inst : compare4 PORT MAP(
		dataa	 => dataa_sig,
		AleB	 => AleB_sig
	);
