count1_inst : count1 PORT MAP(
		clock	 => clock_sig,
		aset	 => aset_sig,
		q	 => q_sig
	);
