compare6_inst : compare6 PORT MAP(
		dataa	 => dataa_sig,
		AeB	 => AeB_sig
	);
