counter1_inst : counter1 PORT MAP(
		clock	 => clock_sig,
		q	 => q_sig
	);
